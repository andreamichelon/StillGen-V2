<?xml version="1.0" encoding="UTF-8"?>
<ColorCorrection id="cc0001">
    <SOPNode>
        <Slope>0.9407 0.9836 0.9794</Slope>
        <Offset>-0.0070 -0.0011 0.0044</Offset>
        <Power>0.9705 1.0210 1.0298</Power>
    </SOPNode>
    <SatNode>
        <Saturation>0.9415</Saturation>
    </SatNode>
</ColorCorrection>